`define NR_REG  32
`define WIDTH   32

`define TLBENTRY    16
