`define NR_REG  32
`define WIDTH   32
