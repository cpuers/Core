module test (
    input x,
    output y
);
    framework u(.x(x), .y(y));
endmodule
