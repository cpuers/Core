module framework (
    input x,
    output y
);
    assign y = x;
endmodule
