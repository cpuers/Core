`ifndef CONFIG_VH
`define CONFIG_VH

`define NR_REG  32
`define WIDTH   32
`define PALEN   32

`define TLBENTRY    16

`endif
